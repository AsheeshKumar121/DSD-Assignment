`timescale 1ns / 1ps

module tb_MUX_8X1(

    );

    reg S0, S1, S2, I0, I1, I2, I3, I4, I5, I6, I7;
    wire Y;

    MUX_8X1 uut (S2, S1, S0, I0, I1, I2, I3, I4, I5, I6, I7, Y);
    initial
    begin
        S0=0; S1=0; S2=0; I0=1; I1=0; I2=0; I3=0; I4=0; I5=0; I6=0; I7=0;
        #10;     
        S0=0; S1=1; S2=0; I0=0; I1=1; I2=0; I3=0; I4=0; I5=0; I6=0; I7=0;
        #10;    
        S0=1; S1=0; S2=0; I0=0; I1=0; I2=1; I3=0; I4=0; I5=0; I6=0; I7=0;
        #10;  
        S0=1; S1=1; S2=0; I0=0; I1=0; I2=0; I3=1; I4=0; I5=0; I6=0; I7=0;
        #10;   
        S0=0; S1=0; S2=1; I0=0; I1=0; I2=0; I3=0; I4=1; I5=0; I6=0; I7=0;
        #10;     
        S0=0; S1=1; S2=1; I0=0; I1=0; I2=0; I3=0; I4=0; I5=1; I6=0; I7=0;
        #10;   
        S0=1; S1=0; S2=1; I0=0; I1=0; I2=0; I3=0; I4=0; I5=0; I6=1; I7=0;
        #10;   
        S0=1; S1=1; S2=1; I0=0; I1=0; I2=0; I3=0; I4=0; I5=0; I6=0; I7=1;
        #10;
        $finish;
    end
endmodule